//Flip Flop de 6 bits
module Flip_D6(input clk, reset,
               input [5:0]d,
               output reg [5:0]q);

  always @(posedge clk, posedge reset) begin
  if (reset) q<=6'b0;
  else       q<=d;
  end
endmodule
//Flip Flop de 3 bits
module Flip_D3(input clk, reset, input [2:0]d, output reg [2:0]q);

    always @ ( posedge clk, posedge reset ) begin
      if (reset) q<=3'b0;
      else       q<=d;
    end
endmodule

//Timer
module Timer(input To, output reg T);

  always @(To)
  if(To == 1) begin
    T = 1;
    #12
    T = 0;
  end
  else
  T = 0;
endmodule

//FSM de Control
module FSM1(input clock, reset, W, A, ES, D,
  input [2:0]E,
  output wire [5:0]SY, SF, S,
  output [3:0]M, YA, AR, F);
//Estados Futuros
  assign SF[5]=(~S[5]&S[4]&S[3]&S[2]&~W&ES&~E[2]&E[1]&E[0])|(S[5]&~S[4]&~S[3]&~S[2]&~W&ES&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&S[3]&S[1]&S[0]&~W&ES&~E[2]&E[1]&E[0])|(~S[5]&S[4]&S[3]&S[2]&~W&A&~D&~E[2]&E[1]&E[0])|
	(S[5]&~S[4]&~S[3]&~S[2]&~W&A&~D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&S[3]&S[2]&A&ES&~D&~E[2]&E[1]&E[0])|
	(S[5]&~S[4]&~S[3]&~S[2]&A&ES&~D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&S[3]&S[1]&S[0]&~W&A&~D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&S[3]&S[1]&S[0]&A&ES&~D&~E[2]&E[1]&E[0]);

  assign SF[4]=(~S[5]&S[4]&~S[3]&~E[2]&E[1]&E[0])|(~S[5]&~S[4]&S[3]&S[2]&~E[2]&E[1]&E[0])|
   (~S[5]&~S[4]&S[3]&S[2]&E[2]&~E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[1]&E[2]&~E[1]&~E[0])|
   (~S[5]&~S[4]&S[3]&S[0]&E[2]&~E[1]&~E[0])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&E[2]&~E[1]&~E[0])|
   (S[5]&~S[4]&~S[3]&~S[2]&W&~A&~E[2]&E[1]&E[0])|(S[5]&~S[4]&~S[3]&~S[2]&W&~ES&~E[2]&E[1]&E[0])|
   (S[5]&~S[4]&~S[3]&~S[2]&~A&~ES&~E[2]&E[1]&E[0])|(S[5]&~S[4]&~S[3]&~S[2]&W&D&~E[2]&E[1]&E[0])|
   (S[5]&~S[4]&~S[3]&~S[2]&~ES&D&~E[2]&E[1]&E[0])|(~S[5]&~S[4]&S[3]&S[2]&~W&A&ES&D&~E[2]&E[1])|
   (~S[5]&~S[4]&S[3]&S[1]&~W&A&ES&D&~E[2]&E[1])|(~S[5]&~S[4]&S[3]&S[0]&~W&A&ES&D&~E[2]&E[1])|
   (~S[5]&~S[4]&S[3]&S[2]&W&A&ES&~D&~E[2]&E[1])|(~S[5]&~S[4]&S[3]&S[1]&W&A&ES&~D&~E[2]&E[1])|
   (~S[5]&~S[4]&S[3]&S[0]&W&A&ES&~D&~E[2]&E[1])|(~S[5]&~S[4]&S[3]&S[2]&~W&~A&ES&~D&~E[2]&E[1])|
   (~S[5]&~S[4]&S[3]&S[1]&~W&~A&ES&~D&~E[2]&E[1])|(~S[5]&~S[4]&S[3]&S[0]&~W&~A&ES&~D&~E[2]&E[1])|
   (~S[5]&~S[4]&S[3]&S[2]&~W&A&~ES&~D&~E[2]&E[1])|(~S[5]&~S[4]&S[3]&S[1]&~W&A&~ES&~D&~E[2]&E[1])|
   (~S[5]&~S[4]&S[3]&S[0]&~W&A&~ES&~D&~E[2]&E[1])|(~S[5]&~S[4]&S[3]&S[2]&~W&A&ES&D&~E[2]&E[0])|
   (~S[5]&~S[4]&S[3]&S[1]&~W&A&ES&D&~E[2]&E[0])|(~S[5]&~S[4]&S[3]&S[0]&~W&A&ES&D&~E[2]&E[0])|
   (~S[5]&~S[4]&S[3]&S[2]&W&A&ES&~D&~E[2]&E[0])|(~S[5]&~S[4]&S[3]&S[1]&W&A&ES&~D&~E[2]&E[0])|
   (~S[5]&~S[4]&S[3]&S[0]&W&A&ES&~D&~E[2]&E[0])|(~S[5]&~S[4]&S[3]&S[2]&~W&~A&ES&~D&~E[2]&E[0])|
   (~S[5]&~S[4]&S[3]&S[1]&~W&~A&ES&~D&~E[2]&E[0])|(~S[5]&~S[4]&S[3]&S[0]&~W&~A&ES&~D&~E[2]&E[0])|
   (~S[5]&~S[4]&S[3]&S[2]&~W&A&~ES&~D&~E[2]&E[0])|(~S[5]&~S[4]&S[3]&S[1]&~W&A&~ES&~D&~E[2]&E[0])|
   (~S[5]&~S[4]&S[3]&S[0]&~W&A&~ES&~D&~E[2]&E[0])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~W&A&ES&D&~E[2]&E[1])|
   (~S[5]&S[4]&~S[3]&~S[2]&~S[1]&W&A&ES&~D&~E[2]&E[1])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~W&~A&ES&~D&~E[2]&E[1])|
   (~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~W&A&~ES&~D&~E[2]&E[1])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~W&A&ES&D&~E[2]&E[0])|
   (~S[5]&S[4]&~S[3]&~S[2]&~S[1]&W&A&ES&~D&~E[2]&E[0])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~W&~A&ES&~D&~E[2]&E[0])|
   (~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~W&A&~ES&~D&~E[2]&E[0])|(~S[5]&~S[4]&S[3]&S[1]&~E[2]&E[1]&E[0])|
   (~S[5]&S[4]&~S[2]&~S[0]&~E[2]&E[1]&E[0])|(~S[5]&S[4]&W&~A&~E[2]&E[1]&E[0])|
   (~S[5]&S[4]&W&~ES&~E[2]&E[1]&E[0])|(~S[5]&S[4]&~A&~ES&~E[2]&E[1]&E[0])|
   (~S[5]&S[4]&W&D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&~ES&D&~E[2]&E[1]&E[0])|
   (~S[5]&S[3]&~S[2]&~S[1]&S[0]&~E[2]&E[1]&E[0]);

assign SF[3]=(~S[5]&~S[4]&~S[3]&~E[2]&~E[1]&E[0])|(~S[5]&~S[4]&W&~A&~E[2]&~E[1]&E[0])|
  (~S[5]&~S[4]&W&~ES&~E[2]&~E[1]&E[0])|(~S[5]&~S[4]&~A&~ES&~E[2]&~E[1]&E[0])|
	(~S[5]&~S[4]&W&D&~E[2]&~E[1]&E[0])|(~S[5]&~S[4]&~A&D&~E[2]&~E[1]&E[0])|
	(~S[5]&~S[4]&~ES&D&~E[2]&~E[1]&E[0])|(~S[5]&~S[4]&S[3]&S[2]&E[2]&~E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[1]&E[2]&~E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[0]&E[2]&~E[1]&~E[0])|
	(~S[5]&~S[4]&~S[2]&~S[1]&~S[0]&~E[2]&~E[1]&E[0])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&E[2]&~E[1]&~E[0])|
	(~S[5]&~S[4]&~S[3]&~W&A&ES&D&~E[2]&~E[1])|(~S[5]&~S[4]&~S[3]&~W&~A&ES&~D&~E[2]&~E[1])|
	(~S[5]&S[4]&S[3]&S[2]&W&~A&~E[2]&E[1]&E[0])|(S[5]&~S[4]&~S[3]&~S[2]&W&~A&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&S[3]&S[2]&W&~ES&~E[2]&E[1]&E[0])|(S[5]&~S[4]&~S[3]&~S[2]&W&~ES&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&S[3]&S[2]&~A&~ES&~E[2]&E[1]&E[0])|(S[5]&~S[4]&~S[3]&~S[2]&~A&~ES&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&S[3]&S[2]&W&D&~E[2]&E[1]&E[0])|(S[5]&~S[4]&~S[3]&~S[2]&W&D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&S[3]&S[2]&~ES&D&~E[2]&E[1]&E[0])|(S[5]&~S[4]&~S[3]&~S[2]&~ES&D&~E[2]&E[1]&E[0])|
	(~S[5]&~S[3]&~S[2]&~S[1]&W&~A&~E[2]&~E[1]&E[0])|(~S[5]&~S[3]&~S[2]&~S[1]&W&~ES&~E[2]&~E[1]&E[0])|
	(~S[5]&~S[3]&~S[2]&~S[1]&~A&~ES&~E[2]&~E[1]&E[0])|(~S[5]&~S[3]&~S[2]&~S[1]&W&D&~E[2]&~E[1]&E[0])|
	(~S[5]&~S[3]&~S[2]&~S[1]&~A&D&~E[2]&~E[1]&E[0])|(~S[5]&~S[3]&~S[2]&~S[1]&~ES&D&~E[2]&~E[1]&E[0])|
	(~S[5]&~S[4]&~W&A&ES&~D&~E[2]&~E[1]&E[0])|(~S[5]&~S[4]&S[3]&S[2]&W&~A&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[1]&W&~A&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[0]&W&~A&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[2]&W&~ES&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[1]&W&~ES&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[0]&W&~ES&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[2]&~A&~ES&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[1]&~A&~ES&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[0]&~A&~ES&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[2]&W&D&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[1]&W&D&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[0]&W&D&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[2]&~A&D&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[1]&~A&D&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[0]&~A&D&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[2]&~ES&D&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[1]&~ES&D&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[0]&~ES&D&~E[2]&E[1]&~E[0])|(~S[5]&S[4]&S[3]&S[1]&S[0]&W&~A&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&~S[3]&S[2]&~W&A&ES&~E[2]&E[1]&E[0])|(~S[5]&S[4]&~S[3]&S[1]&~W&A&ES&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&S[3]&S[1]&S[0]&W&~ES&~E[2]&E[1]&E[0])|(~S[5]&S[4]&S[3]&S[1]&S[0]&~A&~ES&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&S[3]&S[1]&S[0]&W&D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&S[3]&S[1]&S[0]&~ES&D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&~S[3]&S[2]&~W&A&~D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&~S[3]&S[1]&~W&A&~D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&~S[3]&S[2]&~W&ES&~D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&~S[3]&S[1]&~W&ES&~D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&~S[3]&S[2]&A&ES&~D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&~S[3]&S[1]&A&ES&~D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&W&~A&~E[2]&E[1]&~E[0])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&W&~ES&~E[2]&E[1]&~E[0])|
	(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~A&~ES&~E[2]&E[1]&~E[0])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&W&D&~E[2]&E[1]&~E[0])|
	(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~A&D&~E[2]&E[1]&~E[0])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~ES&D&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&~S[2]&~S[1]&~S[0]&~W&A&ES&D&~E[2]&~E[1])|(~S[5]&~S[4]&~S[2]&~S[1]&~S[0]&~W&~A&ES&~D&~E[2]&~E[1])|
	(~S[5]&S[4]&S[3]&~S[2]&~S[1]&~W&A&ES&~E[2]&E[1]&E[0])|(~S[5]&S[4]&S[3]&~S[2]&~S[1]&~W&A&~D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&S[3]&~S[2]&~S[1]&~W&ES&~D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&S[3]&~S[2]&~S[1]&A&ES&~D&~E[2]&E[1]&E[0])|
	(~S[5]&~S[3]&~S[2]&~S[1]&~W&A&ES&~D&~E[2]&~E[1]&E[0])|(~S[5]&~S[4]&S[3]&S[2]&~W&A&ES&~D&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[1]&~W&A&ES&~D&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[0]&~W&A&ES&~D&~E[2]&E[1]&~E[0])|
	(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~W&A&ES&~D&~E[2]&E[1]&~E[0])|(~S[5]&S[4]&~S[2]&S[1]&~S[0]&~W&A&ES&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&~S[2]&S[1]&~S[0]&~W&A&~D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&~S[2]&S[1]&~S[0]&~W&ES&~D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&~S[2]&S[1]&~S[0]&A&ES&~D&~E[2]&E[1]&E[0]);

assign SF[2]=(~S[5]&S[4]&S[3]&S[2]&W&~ES&~E[2]&E[1]&E[0])|(S[5]&~S[4]&~S[3]&~S[2]&W&~ES&~E[2]&E[1]&E[0])|
    (~S[5]&S[4]&~S[3]&S[2]&~A&D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&~S[3]&S[1]&~A&D&~E[2]&E[1]&E[0])|
	(~S[5]&~S[4]&~S[3]&~W&~A&D&~E[2]&~E[1]&~E[0])|(~S[5]&~S[4]&~S[3]&~A&ES&D&~E[2]&~E[1]&~E[0])|
	(~S[5]&~S[4]&~S[3]&~W&A&~D&~E[2]&~E[1]&~E[0])|(~S[5]&~S[4]&~S[3]&A&ES&~D&~E[2]&~E[1]&~E[0])|
	(~S[5]&S[4]&S[3]&S[1]&S[0]&W&~ES&~E[2]&E[1]&E[0])|(~S[5]&S[4]&S[3]&~S[2]&~S[1]&~A&D&~E[2]&E[1]&E[0])|
	(S[5]&~S[4]&~S[3]&~S[2]&W&~A&D&~E[2]&E[1]&E[0])|(S[5]&~S[4]&~S[3]&~S[2]&~A&~ES&D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&S[3]&W&A&~ES&~D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&S[2]&W&A&~ES&~D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&S[1]&W&A&~ES&~D&~E[2]&E[1]&E[0])|(~S[5]&~S[4]&S[3]&S[2]&~W&~A&D&~E[2]&~E[1]&E[0])|
	(~S[5]&~S[4]&S[3]&S[1]&~W&~A&D&~E[2]&~E[1]&E[0])|(~S[5]&~S[4]&S[3]&S[0]&~W&~A&D&~E[2]&~E[1]&E[0])|
	(~S[5]&~S[4]&S[3]&S[2]&~A&ES&D&~E[2]&~E[1]&E[0])|(~S[5]&~S[4]&S[3]&S[1]&~A&ES&D&~E[2]&~E[1]&E[0])|
	(~S[5]&~S[4]&S[3]&S[0]&~A&ES&D&~E[2]&~E[1]&E[0])|(~S[5]&~S[4]&S[3]&S[2]&~W&~A&D&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[1]&~W&~A&D&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[0]&~W&~A&D&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[2]&~A&ES&D&~E[2]&E[1]&~E[0])|(S[5]&~S[4]&S[3]&S[1]&~A&ES&D&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[0]&~A&ES&D&~E[2]&E[1]&~E[0])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~W&~A&D&~E[2]&~E[1]&E[0])|
	(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~A&ES&D&~E[2]&~E[1]&E[0])|(~S[5]&~S[4]&S[3]&S[2]&~W&A&ES&~D&~E[2]&~E[1]&E[0])|
	(~S[5]&~S[4]&S[3]&S[1]&~W&A&ES&~D&~E[2]&~E[1]&E[0])|(~S[5]&~S[4]&S[3]&S[0]&~W&A&ES&~D&~E[2]&~E[1]&E[0])|
	(~S[5]&~S[4]&S[3]&S[2]&W&A&~ES&~D&~E[2]&~E[1]&E[0])|(~S[5]&~S[4]&S[3]&S[1]&W&A&~ES&~D&~E[2]&~E[1]&E[0])|
	(~S[5]&~S[4]&S[3]&S[0]&W&A&~ES&~D&~E[2]&~E[1]&E[0])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~W&~A&D&~E[2]&E[1]&~E[0])|
	(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~A&ES&D&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[2]&~W&A&ES&~D&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[1]&~W&A&ES&~D&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[0]&~W&A&ES&~D&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[2]&W&A&~ES&~D&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[1]&W&A&~ES&~D&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[0]&W&A&~ES&~D&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&~S[2]&~S[1]&~S[0]&~W&~A&D&~E[2]&~E[1]&~E[0])|
	(~S[5]&~S[4]&~S[2]&~S[1]&~S[0]&~A&ES&D&~E[2]&~E[1]&~E[0])|(~S[5]&~S[4]&~S[2]&~S[1]&~S[0]&~W&A&~D&~E[2]&~E[1]&~E[0])|
	(~S[5]&~S[4]&~S[2]&~S[1]&~S[0]&A&ES&~D&~E[2]&~E[1]&~E[0])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~W&A&ES&~D&~E[2]&~E[1]&E[0])|
	(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&W&A&~ES&~D&~E[2]&~E[1]&E[0])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~W&A&ES&~D&~E[2]&E[1]&~E[0])|
	(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&W&A&~ES&~D&~E[2]&E[1]&~E[0])|(~S[5]&S[4]&S[3]&W&~A&D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&S[3]&~A&~ES&D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&~S[2]&S[1]&~S[0]&~A&D&~E[2]&E[1]&E[0]);

assign SF[1]=(~S[5]&~S[4]&S[3]&S[1]&~E[2]&E[1]&E[0])|(~S[5]&~S[4]&S[3]&S[0]&~E[2]&E[1]&E[0])|
    (~S[5]&~S[4]&S[3]&S[2]&E[2]&~E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[1]&E[2]&~E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[0]&E[2]&~E[1]&~E[0])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&~S[3]&A&D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&~S[3]&~A&~D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&E[2]&~E[1]&~E[0])|(~S[5]&~S[4]&~S[3]&A&~D&~E[2]&~E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[2]&W&~A&~ES&~E[2]&E[1])|(~S[5]&~S[4]&S[3]&S[1]&W&~A&~ES&~E[2]&E[1])|
	(~S[5]&~S[4]&S[3]&S[0]&W&~A&~ES&~E[2]&E[1])+(~S[5]&~S[4]&S[3]&S[2]&W&~ES&D&~E[2]&E[1])|
	(~S[5]&~S[4]&S[3]&S[1]&W&~ES&D&~E[2]&E[1])|(~S[5]&~S[4]&S[3]&S[0]&W&~ES&D&~E[2]&E[1])|
	(~S[5]&~S[4]&S[3]&S[2]&W&~A&~ES&~E[2]&E[0])|(~S[5]&~S[4]&S[3]&S[1]&W&~A&~ES&~E[2]&E[0])|
	(~S[5]&~S[4]&S[3]&S[0]&W&~A&~ES&~E[2]&E[0])|(~S[5]&~S[4]&S[3]&S[2]&W&~ES&D&~E[2]&E[0])|
	(~S[5]&~S[4]&S[3]&S[1]&W&~ES&D&~E[2]&E[0])|(~S[5]&~S[4]&S[3]&S[0]&W&~ES&D&~E[2]&E[0])|
	(S[5]&~S[4]&~S[3]&~S[2]&W&ES&~E[2]&E[1]&E[0])|(S[5]&~S[4]&~S[3]&~S[2]&~W&~ES&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&W&~A&~ES&~E[2]&E[1])|(~S[5]&~S[4]&S[3]&S[2]&~W&~A&ES&D&~E[2]&E[1])|
	(~S[5]&~S[4]&S[3]&S[1]&~W&~A&ES&D&~E[2]&E[1])|(~S[5]&~S[4]&S[3]&S[0]&~W&~A&ES&D&~E[2]&E[1])|
	(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&W&~ES&D&~E[2]&E[1])|(~S[5]&~S[4]&S[3]&S[2]&~W&A&ES&~D&~E[2]&E[1])|
	(~S[5]&~S[4]&S[3]&S[1]&~W&A&ES&~D&~E[2]&E[1])|(~S[5]&~S[4]&S[3]&S[0]&~W&A&ES&~D&~E[2]&E[1])|
	(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&W&~A&~ES&~E[2]&E[0])|(~S[5]&~S[4]&S[3]&S[2]&~W&~A&ES&D&~E[2]&E[0])|
	(~S[5]&~S[4]&S[3]&S[1]&~W&~A&ES&D&~E[2]&E[0])|(~S[5]&~S[4]&S[3]&S[0]&~W&~A&ES&D&~E[2]&E[0])|
	(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&W&~ES&D&~E[2]&E[0])|(~S[5]&~S[4]&S[3]&S[2]&~W&A&ES&~D&~E[2]&E[0])|
	(~S[5]&~S[4]&S[3]&S[1]&~W&A&ES&~D&~E[2]&E[0])|(~S[5]&~S[4]&S[3]&S[0]&~W&A&ES&~D&~E[2]&E[0])|
	(~S[5]&~S[4]&~S[3]&W&~A&~ES&D&~E[2]&~E[1]&~E[0])|(~S[5]&~S[4]&~S[2]&~S[1]&~S[0]&A&~D&~E[2]&~E[1]&~E[0])|
	(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~W&~A&ES&D&~E[2]&E[1])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~W&A&ES&~D&~E[2]&E[1])|
	(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~W&~A&ES&D&~E[2]&E[0])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~W&A&ES&~D&~E[2]&E[0])|
	(~S[5]&~S[4]&~S[2]&~S[1]&~S[0]&W&~A&~ES&D&~E[2]&~E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[2]&~E[2]&E[1]&E[0])|
	(~S[5]&S[3]&S[2]&~W&~ES&~E[2]&E[1]&E[0])|(~S[5]&S[4]&~S[3]&~W&D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&W&ES&D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&A&ES&D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&~A&ES&~D&~E[2]&E[1]&E[0])|(~S[5]&S[3]&S[1]&S[0]&~W&~ES&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&~S[2]&~S[1]&~W&D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&~S[2]&~S[0]&~W&D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&~S[2]&~S[1]&A&D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&~S[2]&~S[0]&A&D&~E[2]&E[1]&E[0])|
	(~S[5]&S[3]&S[2]&W&A&~D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&~S[2]&~S[1]&~A&~D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&~S[2]&~S[0]&~A&~D&~E[2]&E[1]&E[0])|(S[5]&~S[4]&~S[3]&~S[2]&A&ES&D&~E[2]&E[1]&E[0])|
	(~S[5]&S[3]&S[1]&S[0]&W&A&~D&~E[2]&E[1]&E[0])|(S[5]&~S[4]&~S[3]&~S[2]&~A&ES&~D&~E[2]&E[1]&E[0])|
	(S[5]&~S[4]&~S[3]&~S[2]&A&~ES&~D&~E[2]&E[1]&E[0]);

assign SF[0]=(~S[5]&~S[4]&S[3]&S[2]&E[2]&~E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[1]&E[2]&~E[1]&~E[0])|
    (~S[5]&~S[4]&S[3]&S[0]&E[2]&~E[1]&~E[0])|(~S[5]&~S[4]&~S[3]&W&A&~ES&~E[2]&~E[1])|
	(~S[5]&~S[4]&~S[3]&W&A&~D&~E[2]&~E[1])|(~S[5]&~S[4]&~S[3]&W&~ES&~D&~E[2]&~E[1])|
	(~S[5]&~S[4]&~S[3]&A&~ES&~D&~E[2]&~E[1])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&E[2]&~E[1]&~E[0])|
	(~S[5]&~S[4]&~S[3]&~W&~A&ES&D&~E[2]&~E[1])|(~S[5]&~S[4]&~S[2]&~S[1]&~S[0]&W&A&~ES&~E[2]&~E[1])|
	(~S[5]&~S[4]&~S[2]&~S[1]&~S[0]&W&A&~D&~E[2]&~E[1])|(~S[5]&~S[4]&~S[2]&~S[1]&~S[0]&W&~ES&~D&~E[2]&~E[1])|
	(~S[5]&~S[4]&~S[2]&~S[1]&~S[0]&A&~ES&~D&~E[2]&~E[1])|(~S[5]&S[4]&~S[3]&S[2]&W&A&~ES&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&~S[3]&S[1]&W&A&~ES&~E[2]&E[1]&E[0])|(~S[5]&S[4]&~S[3]&S[2]&W&A&~D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&~S[3]&S[1]&W&A&~D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&~S[3]&S[2]&W&~ES&~D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&~S[3]&S[1]&W&~ES&~D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&~S[3]&S[2]&A&~ES&~D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&~S[3]&S[1]&A&~ES&~D&~E[2]&E[1]&E[0])|(~S[5]&~S[4]&~S[2]&~S[1]&~S[0]&~W&~A&ES&D&~E[2]&~E[1])|
	(~S[5]&S[4]&S[3]&~S[2]&~S[1]&W&A&~ES&~E[2]&E[1]&E[0])|(~S[5]&S[4]&~S[3]&S[2]&~W&~A&ES&D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&~S[3]&S[1]&~W&~A&ES&D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&S[3]&~S[2]&~S[1]&W&A&~D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&S[3]&~S[2]&~S[1]&W&~ES&~D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&S[3]&~S[2]&~S[1]&A&~ES&~D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&S[3]&~S[2]&~S[1]&~W&~A&ES&D&~E[2]&E[1]&E[0])|(~S[5]&~S[4]&W&~A&ES&~E[2]&~E[1]&E[0])|
	(~S[5]&~S[4]&~W&~A&~ES&~E[2]&~E[1]&E[0])|(~S[5]&~S[4]&A&ES&D&~E[2]&~E[1]&E[0])|
	(~S[5]&~S[4]&~W&~ES&D&~E[2]&~E[1]&E[0])|(~S[5]&~S[4]&~A&~ES&D&~E[2]&~E[1]&E[0])|
	(~S[5]&~S[4]&~W&ES&~D&~E[2]&~E[1]&E[0])|(~S[5]&S[4]&S[3]&S[2]&W&~A&ES&~E[2]&E[1]&E[0])|
	(S[5]&~S[4]&~S[3]&~S[2]&W&~A&ES&~E[2]&E[1]&E[0])|(~S[5]&S[4]&S[3]&S[2]&~W&~A&~ES&~E[2]&E[1]&E[0])|
	(S[5]&~S[4]&~S[3]&~S[2]&~W&~A&~ES&~E[2]&E[1]&E[0])|(~S[5]&S[4]&S[3]&S[2]&A&ES&D&~E[2]&E[1]&E[0])|
	(S[5]&~S[4]&~S[3]&~S[2]&A&ES&D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&S[3]&S[2]&~W&~ES&D&~E[2]&E[1]&E[0])|
	(S[5]&~S[4]&~S[3]&~S[2]&~W&~ES&D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&S[3]&S[2]&~A&~ES&D&~E[2]&E[1]&E[0])|
	(S[5]&~S[4]&~S[3]&~S[2]&~A&~ES&D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&S[3]&S[2]&~W&ES&~D&~E[2]&E[1]&E[0])|
	(S[5]&~S[4]&~S[3]&~S[2]&~W&ES&~D&~E[2]&E[1]&E[0])|(~S[5]&~S[3]&~S[2]&~S[1]&W&~A&ES&~E[2]&~E[1]&E[0])|
	(~S[5]&~S[3]&~S[2]&~S[1]&~W&~A&~ES&~E[2]&~E[1]&E[0])|(~S[5]&~S[3]&~S[2]&~S[1]&A&ES&D&~E[2]&~E[1]&E[0])|
	(~S[5]&~S[3]&~S[2]&~S[1]&~W&~ES&D&~E[2]&~E[1]&E[0])|(~S[5]&~S[3]&~S[2]&~S[1]&~A&~ES&D&~E[2]&~E[1]&E[0])|
	(~S[5]&~S[3]&~S[2]&~S[1]&~W&ES&~D&~E[2]&~E[1]&E[0])|(~S[5]&~S[4]&S[3]&S[2]&W&~A&ES&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[1]&W&~A&ES&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[0]&W&~A&ES&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[2]&~W&~A&~ES&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[1]&~W&~A&~ES&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[0]&~W&~A&~ES&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[2]&A&ES&D&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[1]&A&ES&D&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[0]&A&ES&D&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[2]&~W&~ES&D&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[1]&~W&~ES&D&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[0]&~W&~ES&D&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[2]&~A&~ES&D&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[1]&~A&~ES&D&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[0]&~A&~ES&D&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[2]&~W&ES&~D&~E[2]&E[1]&~E[0])|(~S[5]&~S[4]&S[3]&S[1]&~W&ES&~D&~E[2]&E[1]&~E[0])|
	(~S[5]&~S[4]&S[3]&S[0]&~W&ES&~D&~E[2]&E[1]&~E[0])|(~S[5]&S[4]&S[3]&S[1]&S[0]&W&~A&ES&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&~S[2]&S[1]&~S[0]&W&A&~ES&~E[2]&E[1]&E[0])|(~S[5]&S[4]&S[3]&S[1]&S[0]&~W&~A&~ES&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&S[3]&S[1]&S[0]&A&ES&D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&S[3]&S[1]&S[0]&~W&~ES&D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&S[3]&S[1]&S[0]&~A&~ES&D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&~S[2]&S[1]&~S[0]&W&A&~D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&S[3]&S[1]&S[0]&~W&ES&~D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&~S[2]&S[1]&~S[0]&W&~ES&~D&~E[2]&E[1]&E[0])|
	(~S[5]&S[4]&~S[2]&S[1]&~S[0]&A&~ES&~D&~E[2]&E[1]&E[0])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&W&~A&ES&~E[2]&E[1]&~E[0])|
	(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~W&~A&~ES&~E[2]&E[1]&~E[0])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&A&ES&D&~E[2]&E[1]&~E[0])|
	(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~W&~ES&D&~E[2]&E[1]&~E[0])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~A&~ES&D&~E[2]&E[1]&~E[0])|
	(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~W&ES&~D&~E[2]&E[1]&~E[0])|(~S[5]&S[4]&~S[2]&S[1]&~S[0]&~W&~A&ES&D&~E[2]&E[1]&E[0]);
//Salidas
assign SY[5]=S[5];
assign SY[4]=S[4];
assign SY[3]=S[3];
assign SY[2]=S[2];
assign SY[1]=S[1];
assign SY[0]=S[0];
assign M[3]=~S[5]&~S[4]&S[3]&~S[2]&~S[1]&~S[0];
assign M[2]=~S[5]&~S[4]&~S[3]&S[2];
assign M[1]=~S[5]&~S[4]&~S[3]&S[1];
assign M[0]=~S[5]&~S[4]&~S[3]&S[0];
assign YA[3]=~S[5]&S[4]&~S[3]&~S[2]&~S[1]&S[0];
assign YA[2]=(~S[5]&~S[4]&S[3]&S[2]&S[1])|(~S[5]&~S[4]&S[3]&S[2]&S[0])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~S[0]);
assign YA[1]=(~S[5]&~S[4]&S[3]&S[1]&S[0])|(~S[5]&~S[4]&S[3]&S[2]&~S[1]&~S[0])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~S[0]);
assign YA[0]=(~S[5]&~S[4]&S[3]&S[2]&~S[0])|(~S[5]&~S[4]&S[3]&S[1]&~S[0])|(~S[5]&S[4]&~S[3]&~S[2]&~S[1]&~S[0]);
assign F[3]=~S[5]&S[4]&S[3]&~S[2]&S[1]&~S[0];
assign F[2]=(~S[5]&S[4]&~S[3]&S[2]&S[1])|(~S[5]&S[4]&S[3]&~S[2]&~S[1]);
assign F[1]=(~S[5]&S[4]&~S[3]&S[2]&~S[1])|(~S[5]&S[4]&S[3]&~S[2]&~S[1]);
assign F[0]=(~S[5]&S[4]&~S[3]&S[2]&S[0])|(~S[5]&S[4]&~S[3]&S[1]&S[0])|(~S[5]&S[4]&S[3]&~S[2]&~S[1]&S[0]);
assign AR[3]=S[5]&~S[4]&~S[3]&~S[2]&S[1]&S[0];
assign AR[2]=(S[5]&~S[4]&~S[3]&~S[2]&~S[1])|(S[5]&~S[4]&~S[3]&~S[2]&~S[0])|(~S[5]&S[4]&S[3]&S[2]&S[1]&S[0]);
assign AR[1]=(~S[5]&S[4]&S[3]&S[2]&~S[1]&S[0])|(S[5]&~S[4]&~S[3]&~S[2]&~S[1]&S[0])|(~S[5]&S[4]&S[3]&S[2]&S[1]&~S[0])|(S[5]&~S[4]&~S[3]&~S[2]&S[1]&~S[0]);
assign AR[0]=(~S[5]&S[4]&S[3]&S[2]&~S[0])|(S[5]&~S[4]&~S[3]&~S[2]&~S[0]);

Flip_D6 U6(.clk(clock), .reset(reset), .d(SF), .q(S));

endmodule
//FMS de Estados
module FSM2(input clock, reset, SLT, R, T,
  output To,
  output wire [2:0] SY,SF, S);
//Estados Futuros
assign SF[2] = (S[2]&~S[1]&~S[0]&T)|(~S[2]&S[1]&~S[0]&~SLT&T&R);
assign SF[1] = (~S[2]&~S[1]&S[0])|(~S[2]&S[0]&T)|(~S[2]&S[1]&SLT&T)|(~S[2]&S[1]&T&~R);
assign SF[0] = (~S[2]&S[1]&S[0]&T)|(~S[2]&S[1]&SLT&T)|(~S[2]&~S[1]&~S[0]&SLT&~T);
//Salidas
assign SY[2]=S[2];
assign SY[1]=S[1];
assign SY[0]=S[0];
assign To = (~S[2]&~S[1]&S[0])|(~S[2]&S[1]&~S[0])|(~S[2]&S[1]&S[0])|(S[2]&~S[1]&~S[0]);
Flip_D3 U5(.clk(clock), .reset(reset), .d(SF), .q(S));
endmodule
module Proyecto1(input wire clock1, reset1, W, A, ES, D, SLT2, R2, T,
              output wire [3:0]M, YA, AR, F);
              wire g, TOS;
              wire [3:0]C3, C4, C5, C6, C7;
              wire [2:0]C2, C8, C9;
              wire [5:0]C1, C10, C11;

              FSM2 U1(.clock(clock1), .reset(reset1), .SLT(SLT2),  .R(R2),  .T(T), .To(TOS), .SY(C2), .SF(C8), .S(C9));
              Timer U2(.To(TOS), .T(g));
              FSM1 U3(.clock(clock1), .reset(reset1), .W(W), .A(A), .ES(ES), .D(D), .E(C2), .SY(C1), .SF(C10), .S(C11), .M(C3), .YA(C4), .AR(C5), .F(C6));
endmodule
